library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

-- Please start to write a entity block ! --



-- End of  a entity block.  --

architecture logic of adder is
begin
	sum <= a + b;
end;